// HMTH (c)

module XAFifo #(parameter DEPTH = 4, DW = 8, W_SYNC_N = 2, R_SYNC_N = 2) (
    input  logic rclk
  , input  logic rrstn

  , input  logic re
  , output logic empty_n

  , input  logic wclk
  , input  logic wrstn

  , input  logic we
  , output logic full_n

	, input  logic [DW-1:0] din
	, output logic [DW-1:0] dout
);

logic                       we_ok;
logic [$clog2(DEPTH) : 0]   a_g_wptr;
logic [$clog2(DEPTH) : 0]   a_g_rptr;

logic [$clog2(DEPTH)-1 : 0] rptr;
logic [$clog2(DEPTH)-1 : 0] wptr;

XAFifoWCtrl #(.DEPTH(DEPTH), .SYNC_N(W_SYNC_N))
	WCtrl (.clk(wclk), .rstn(wrstn), .we(we), .full_n(full_n), .a_g_rptr(a_g_rptr), .a_g_wptr(a_g_wptr), .we_ok(we_ok), .wptr(wptr));

XAFifoRCtrl #(.DEPTH(DEPTH), .SYNC_N(R_SYNC_N))
	RCtrl (.clk(rclk), .rstn(rrstn), .re(re), .empty_n(empty_n), .a_g_rptr(a_g_rptr), .a_g_wptr(a_g_wptr), .rptr(rptr));

XMem #(.DW(DW), .DEPTH(DEPTH))
	Mem (.clk(wclk), .we(we_ok), .waddr(wptr), .raddr(rptr), .d(din), .q(dout));

endmodule

module XAFifoWCtrl #(parameter DEPTH = 4, SYNC_N = 2) (
    input  logic clk
  , input  logic rstn

  , input  logic we
  , output logic full_n

  , input  logic [$clog2(DEPTH) : 0]   a_g_rptr
  , output logic                       we_ok
  , output logic [$clog2(DEPTH)-1 : 0] wptr
  , output logic [$clog2(DEPTH) : 0]   a_g_wptr
);

localparam AW = $clog2(DEPTH);

logic [AW:0] synced_g_rptr;
logic [AW:0] nxt_bin_cnt, bin_cnt, nxt_g_wptr;

XMultiBitSyncer #(.DW(AW+1), .N(SYNC_N)) rptr_syncer (.clk(clk), .rstn(rstn), .d(a_g_rptr), .q(synced_g_rptr));

`ifndef SELECT_SRSTn 
always @(posedge clk, negedge rstn) begin
`else
always @(posedge clk) begin
`endif
  if (~rstn) begin
    bin_cnt                        <= {(AW+1){1'b0}};
    a_g_wptr                       <= {(AW+1){1'b0}};
    full_n                         <= 1'b1;
  end else begin
    bin_cnt                        <= nxt_bin_cnt;
    a_g_wptr                       <= nxt_g_wptr;
    full_n                         <= (nxt_g_wptr [AW] != synced_g_rptr [AW]) && (nxt_g_wptr [AW-1] == ~synced_g_rptr [AW-1]) && (nxt_g_wptr [AW-2:0] == synced_g_rptr [AW-2:0]) ? 1'b0 : 1'b1;
  end
end

assign wptr  = bin_cnt [AW-1:0];
assign we_ok = we & full_n;

assign nxt_bin_cnt = we_ok ? bin_cnt + 1'b1 : bin_cnt;
assign nxt_g_wptr  = (nxt_bin_cnt >> 1) ^ nxt_bin_cnt;

endmodule

module XAFifoRCtrl #(parameter DEPTH = 4, SYNC_N = 2) (
    input  logic clk
  , input  logic rstn

  , input  logic re
  , output logic empty_n

  , input  logic [$clog2(DEPTH) : 0]   a_g_wptr
  , output logic [$clog2(DEPTH)-1 : 0] rptr
  , output logic [$clog2(DEPTH) : 0]   a_g_rptr
);

localparam AW = $clog2(DEPTH);

logic        re_ok;
logic [AW:0] synced_g_wptr;
logic [AW:0] nxt_bin_cnt, bin_cnt, nxt_g_rptr;

XMultiBitSyncer #(.DW(AW+1), .N(SYNC_N)) wptr_syncer (.clk(clk), .rstn(rstn), .d(a_g_wptr), .q(synced_g_wptr));

`ifndef SELECT_SRSTn 
always @(posedge clk, negedge rstn) begin
`else
always @(posedge clk) begin
`endif
  if (~rstn) begin
    bin_cnt                        <= {(AW+1){1'b0}};
    a_g_rptr                       <= {(AW+1){1'b0}};
    empty_n                        <= 1'b0;
  end else begin
    bin_cnt                        <= nxt_bin_cnt;
    a_g_rptr                       <= nxt_g_rptr;
    empty_n                        <= synced_g_wptr == nxt_g_rptr ? 1'b0 : 1'b1;
  end
end

assign rptr  = bin_cnt [AW-1:0];
assign re_ok = re & empty_n;

assign nxt_bin_cnt = re_ok ? bin_cnt + 1'b1 : bin_cnt;
assign nxt_g_rptr  = (nxt_bin_cnt >> 1) ^ nxt_bin_cnt;

endmodule
// EOF
